library ex4_lib1;
use ex4_lib1.lib1;

package ex4 is

    constant ex4_const: integer := lib1.c;

end package ex4;
