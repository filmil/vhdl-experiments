-- The library here is ex4_lib1.

package lib1 is
    
   -- This is ex4_lib1.lib1.c
   constant c: integer := 1; 
    
end package lib1;
